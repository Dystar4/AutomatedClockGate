

module spm
(
  clk,
  rst,
  x,
  y,
  p
);

  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire \$genblock$spm.v:14$10[10].csa.clk ;
  wire \$genblock$spm.v:14$10[10].csa.hsum2 ;
  wire \$genblock$spm.v:14$10[10].csa.rst ;
  wire \$genblock$spm.v:14$10[10].csa.sc ;
  wire \$genblock$spm.v:14$10[10].csa.sum ;
  wire \$genblock$spm.v:14$10[10].csa.y ;
  wire \$genblock$spm.v:14$11[11].csa.clk ;
  wire \$genblock$spm.v:14$11[11].csa.hsum2 ;
  wire \$genblock$spm.v:14$11[11].csa.rst ;
  wire \$genblock$spm.v:14$11[11].csa.sc ;
  wire \$genblock$spm.v:14$11[11].csa.sum ;
  wire \$genblock$spm.v:14$11[11].csa.y ;
  wire \$genblock$spm.v:14$12[12].csa.clk ;
  wire \$genblock$spm.v:14$12[12].csa.hsum2 ;
  wire \$genblock$spm.v:14$12[12].csa.rst ;
  wire \$genblock$spm.v:14$12[12].csa.sc ;
  wire \$genblock$spm.v:14$12[12].csa.sum ;
  wire \$genblock$spm.v:14$12[12].csa.y ;
  wire \$genblock$spm.v:14$13[13].csa.clk ;
  wire \$genblock$spm.v:14$13[13].csa.hsum2 ;
  wire \$genblock$spm.v:14$13[13].csa.rst ;
  wire \$genblock$spm.v:14$13[13].csa.sc ;
  wire \$genblock$spm.v:14$13[13].csa.sum ;
  wire \$genblock$spm.v:14$13[13].csa.y ;
  wire \$genblock$spm.v:14$14[14].csa.clk ;
  wire \$genblock$spm.v:14$14[14].csa.hsum2 ;
  wire \$genblock$spm.v:14$14[14].csa.rst ;
  wire \$genblock$spm.v:14$14[14].csa.sc ;
  wire \$genblock$spm.v:14$14[14].csa.sum ;
  wire \$genblock$spm.v:14$14[14].csa.y ;
  wire \$genblock$spm.v:14$15[15].csa.clk ;
  wire \$genblock$spm.v:14$15[15].csa.hsum2 ;
  wire \$genblock$spm.v:14$15[15].csa.rst ;
  wire \$genblock$spm.v:14$15[15].csa.sc ;
  wire \$genblock$spm.v:14$15[15].csa.sum ;
  wire \$genblock$spm.v:14$15[15].csa.y ;
  wire \$genblock$spm.v:14$16[16].csa.clk ;
  wire \$genblock$spm.v:14$16[16].csa.hsum2 ;
  wire \$genblock$spm.v:14$16[16].csa.rst ;
  wire \$genblock$spm.v:14$16[16].csa.sc ;
  wire \$genblock$spm.v:14$16[16].csa.sum ;
  wire \$genblock$spm.v:14$16[16].csa.y ;
  wire \$genblock$spm.v:14$17[17].csa.clk ;
  wire \$genblock$spm.v:14$17[17].csa.hsum2 ;
  wire \$genblock$spm.v:14$17[17].csa.rst ;
  wire \$genblock$spm.v:14$17[17].csa.sc ;
  wire \$genblock$spm.v:14$17[17].csa.sum ;
  wire \$genblock$spm.v:14$17[17].csa.y ;
  wire \$genblock$spm.v:14$18[18].csa.clk ;
  wire \$genblock$spm.v:14$18[18].csa.hsum2 ;
  wire \$genblock$spm.v:14$18[18].csa.rst ;
  wire \$genblock$spm.v:14$18[18].csa.sc ;
  wire \$genblock$spm.v:14$18[18].csa.sum ;
  wire \$genblock$spm.v:14$18[18].csa.y ;
  wire \$genblock$spm.v:14$19[19].csa.clk ;
  wire \$genblock$spm.v:14$19[19].csa.hsum2 ;
  wire \$genblock$spm.v:14$19[19].csa.rst ;
  wire \$genblock$spm.v:14$19[19].csa.sc ;
  wire \$genblock$spm.v:14$19[19].csa.sum ;
  wire \$genblock$spm.v:14$19[19].csa.y ;
  wire \$genblock$spm.v:14$1[1].csa.clk ;
  wire \$genblock$spm.v:14$1[1].csa.hsum2 ;
  wire \$genblock$spm.v:14$1[1].csa.rst ;
  wire \$genblock$spm.v:14$1[1].csa.sc ;
  wire \$genblock$spm.v:14$1[1].csa.sum ;
  wire \$genblock$spm.v:14$1[1].csa.y ;
  wire \$genblock$spm.v:14$20[20].csa.clk ;
  wire \$genblock$spm.v:14$20[20].csa.hsum2 ;
  wire \$genblock$spm.v:14$20[20].csa.rst ;
  wire \$genblock$spm.v:14$20[20].csa.sc ;
  wire \$genblock$spm.v:14$20[20].csa.sum ;
  wire \$genblock$spm.v:14$20[20].csa.y ;
  wire \$genblock$spm.v:14$21[21].csa.clk ;
  wire \$genblock$spm.v:14$21[21].csa.hsum2 ;
  wire \$genblock$spm.v:14$21[21].csa.rst ;
  wire \$genblock$spm.v:14$21[21].csa.sc ;
  wire \$genblock$spm.v:14$21[21].csa.sum ;
  wire \$genblock$spm.v:14$21[21].csa.y ;
  wire \$genblock$spm.v:14$22[22].csa.clk ;
  wire \$genblock$spm.v:14$22[22].csa.hsum2 ;
  wire \$genblock$spm.v:14$22[22].csa.rst ;
  wire \$genblock$spm.v:14$22[22].csa.sc ;
  wire \$genblock$spm.v:14$22[22].csa.sum ;
  wire \$genblock$spm.v:14$22[22].csa.y ;
  wire \$genblock$spm.v:14$23[23].csa.clk ;
  wire \$genblock$spm.v:14$23[23].csa.hsum2 ;
  wire \$genblock$spm.v:14$23[23].csa.rst ;
  wire \$genblock$spm.v:14$23[23].csa.sc ;
  wire \$genblock$spm.v:14$23[23].csa.sum ;
  wire \$genblock$spm.v:14$23[23].csa.y ;
  wire \$genblock$spm.v:14$24[24].csa.clk ;
  wire \$genblock$spm.v:14$24[24].csa.hsum2 ;
  wire \$genblock$spm.v:14$24[24].csa.rst ;
  wire \$genblock$spm.v:14$24[24].csa.sc ;
  wire \$genblock$spm.v:14$24[24].csa.sum ;
  wire \$genblock$spm.v:14$24[24].csa.y ;
  wire \$genblock$spm.v:14$25[25].csa.clk ;
  wire \$genblock$spm.v:14$25[25].csa.hsum2 ;
  wire \$genblock$spm.v:14$25[25].csa.rst ;
  wire \$genblock$spm.v:14$25[25].csa.sc ;
  wire \$genblock$spm.v:14$25[25].csa.sum ;
  wire \$genblock$spm.v:14$25[25].csa.y ;
  wire \$genblock$spm.v:14$26[26].csa.clk ;
  wire \$genblock$spm.v:14$26[26].csa.hsum2 ;
  wire \$genblock$spm.v:14$26[26].csa.rst ;
  wire \$genblock$spm.v:14$26[26].csa.sc ;
  wire \$genblock$spm.v:14$26[26].csa.sum ;
  wire \$genblock$spm.v:14$26[26].csa.y ;
  wire \$genblock$spm.v:14$27[27].csa.clk ;
  wire \$genblock$spm.v:14$27[27].csa.hsum2 ;
  wire \$genblock$spm.v:14$27[27].csa.rst ;
  wire \$genblock$spm.v:14$27[27].csa.sc ;
  wire \$genblock$spm.v:14$27[27].csa.sum ;
  wire \$genblock$spm.v:14$27[27].csa.y ;
  wire \$genblock$spm.v:14$28[28].csa.clk ;
  wire \$genblock$spm.v:14$28[28].csa.hsum2 ;
  wire \$genblock$spm.v:14$28[28].csa.rst ;
  wire \$genblock$spm.v:14$28[28].csa.sc ;
  wire \$genblock$spm.v:14$28[28].csa.sum ;
  wire \$genblock$spm.v:14$28[28].csa.y ;
  wire \$genblock$spm.v:14$29[29].csa.clk ;
  wire \$genblock$spm.v:14$29[29].csa.hsum2 ;
  wire \$genblock$spm.v:14$29[29].csa.rst ;
  wire \$genblock$spm.v:14$29[29].csa.sc ;
  wire \$genblock$spm.v:14$29[29].csa.sum ;
  wire \$genblock$spm.v:14$29[29].csa.y ;
  wire \$genblock$spm.v:14$2[2].csa.clk ;
  wire \$genblock$spm.v:14$2[2].csa.hsum2 ;
  wire \$genblock$spm.v:14$2[2].csa.rst ;
  wire \$genblock$spm.v:14$2[2].csa.sc ;
  wire \$genblock$spm.v:14$2[2].csa.sum ;
  wire \$genblock$spm.v:14$2[2].csa.y ;
  wire \$genblock$spm.v:14$30[30].csa.clk ;
  wire \$genblock$spm.v:14$30[30].csa.hsum2 ;
  wire \$genblock$spm.v:14$30[30].csa.rst ;
  wire \$genblock$spm.v:14$30[30].csa.sc ;
  wire \$genblock$spm.v:14$30[30].csa.sum ;
  wire \$genblock$spm.v:14$30[30].csa.y ;
  wire \$genblock$spm.v:14$3[3].csa.clk ;
  wire \$genblock$spm.v:14$3[3].csa.hsum2 ;
  wire \$genblock$spm.v:14$3[3].csa.rst ;
  wire \$genblock$spm.v:14$3[3].csa.sc ;
  wire \$genblock$spm.v:14$3[3].csa.sum ;
  wire \$genblock$spm.v:14$3[3].csa.y ;
  wire \$genblock$spm.v:14$4[4].csa.clk ;
  wire \$genblock$spm.v:14$4[4].csa.hsum2 ;
  wire \$genblock$spm.v:14$4[4].csa.rst ;
  wire \$genblock$spm.v:14$4[4].csa.sc ;
  wire \$genblock$spm.v:14$4[4].csa.sum ;
  wire \$genblock$spm.v:14$4[4].csa.y ;
  wire \$genblock$spm.v:14$5[5].csa.clk ;
  wire \$genblock$spm.v:14$5[5].csa.hsum2 ;
  wire \$genblock$spm.v:14$5[5].csa.rst ;
  wire \$genblock$spm.v:14$5[5].csa.sc ;
  wire \$genblock$spm.v:14$5[5].csa.sum ;
  wire \$genblock$spm.v:14$5[5].csa.y ;
  wire \$genblock$spm.v:14$6[6].csa.clk ;
  wire \$genblock$spm.v:14$6[6].csa.hsum2 ;
  wire \$genblock$spm.v:14$6[6].csa.rst ;
  wire \$genblock$spm.v:14$6[6].csa.sc ;
  wire \$genblock$spm.v:14$6[6].csa.sum ;
  wire \$genblock$spm.v:14$6[6].csa.y ;
  wire \$genblock$spm.v:14$7[7].csa.clk ;
  wire \$genblock$spm.v:14$7[7].csa.hsum2 ;
  wire \$genblock$spm.v:14$7[7].csa.rst ;
  wire \$genblock$spm.v:14$7[7].csa.sc ;
  wire \$genblock$spm.v:14$7[7].csa.sum ;
  wire \$genblock$spm.v:14$7[7].csa.y ;
  wire \$genblock$spm.v:14$8[8].csa.clk ;
  wire \$genblock$spm.v:14$8[8].csa.hsum2 ;
  wire \$genblock$spm.v:14$8[8].csa.rst ;
  wire \$genblock$spm.v:14$8[8].csa.sc ;
  wire \$genblock$spm.v:14$8[8].csa.sum ;
  wire \$genblock$spm.v:14$8[8].csa.y ;
  wire \$genblock$spm.v:14$9[9].csa.clk ;
  wire \$genblock$spm.v:14$9[9].csa.hsum2 ;
  wire \$genblock$spm.v:14$9[9].csa.rst ;
  wire \$genblock$spm.v:14$9[9].csa.sc ;
  wire \$genblock$spm.v:14$9[9].csa.sum ;
  wire \$genblock$spm.v:14$9[9].csa.y ;
  input clk;
  wire \csa0.clk ;
  wire \csa0.hsum2 ;
  wire \csa0.rst ;
  wire \csa0.sc ;
  wire \csa0.sum ;
  wire \csa0.y ;
  output p;
  wire [31:1] pp;
  input rst;
  wire \tcmp.clk ;
  wire \tcmp.rst ;
  wire \tcmp.s ;
  wire \tcmp.z ;
  input [31:0] x;
  input y;

  sky130_fd_sc_hd__inv_1
  _223_
  (
    .A(rst),
    .Y(_000_)
  );


  sky130_fd_sc_hd__nand2_1
  _224_
  (
    .A(y),
    .B(x[10]),
    .Y(_045_)
  );


  sky130_fd_sc_hd__nand2_1
  _225_
  (
    .A(\$genblock$spm.v:14$10[10].csa.sc ),
    .B(\$genblock$spm.v:14$11[11].csa.sum ),
    .Y(_046_)
  );


  sky130_fd_sc_hd__nor2_1
  _226_
  (
    .A(\$genblock$spm.v:14$10[10].csa.sc ),
    .B(\$genblock$spm.v:14$11[11].csa.sum ),
    .Y(_047_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _227_
  (
    .A(_046_),
    .SLEEP(_047_),
    .X(_048_)
  );


  sky130_fd_sc_hd__xnor2_1
  _228_
  (
    .A(_045_),
    .B(_048_),
    .Y(\$genblock$spm.v:14$10[10].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _229_
  (
    .A1(_045_),
    .A2(_047_),
    .B1(_046_),
    .Y(_214_)
  );


  sky130_fd_sc_hd__inv_1
  _230_
  (
    .A(rst),
    .Y(_215_)
  );


  sky130_fd_sc_hd__nand2_1
  _231_
  (
    .A(y),
    .B(x[11]),
    .Y(_050_)
  );


  sky130_fd_sc_hd__nand2_1
  _232_
  (
    .A(\$genblock$spm.v:14$11[11].csa.sc ),
    .B(\$genblock$spm.v:14$12[12].csa.sum ),
    .Y(_052_)
  );


  sky130_fd_sc_hd__nor2_1
  _233_
  (
    .A(\$genblock$spm.v:14$11[11].csa.sc ),
    .B(\$genblock$spm.v:14$12[12].csa.sum ),
    .Y(_054_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _234_
  (
    .A(_052_),
    .SLEEP(_054_),
    .X(_055_)
  );


  sky130_fd_sc_hd__xnor2_1
  _235_
  (
    .A(_050_),
    .B(_055_),
    .Y(\$genblock$spm.v:14$11[11].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _236_
  (
    .A1(_050_),
    .A2(_054_),
    .B1(_052_),
    .Y(_216_)
  );


  sky130_fd_sc_hd__inv_1
  _237_
  (
    .A(rst),
    .Y(_217_)
  );


  sky130_fd_sc_hd__inv_1
  _238_
  (
    .A(rst),
    .Y(_218_)
  );


  sky130_fd_sc_hd__nand2_1
  _239_
  (
    .A(y),
    .B(x[12]),
    .Y(_056_)
  );


  sky130_fd_sc_hd__nand2_1
  _240_
  (
    .A(\$genblock$spm.v:14$12[12].csa.sc ),
    .B(\$genblock$spm.v:14$13[13].csa.sum ),
    .Y(_058_)
  );


  sky130_fd_sc_hd__nor2_1
  _241_
  (
    .A(\$genblock$spm.v:14$12[12].csa.sc ),
    .B(\$genblock$spm.v:14$13[13].csa.sum ),
    .Y(_060_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _242_
  (
    .A(_058_),
    .SLEEP(_060_),
    .X(_062_)
  );


  sky130_fd_sc_hd__xnor2_1
  _243_
  (
    .A(_056_),
    .B(_062_),
    .Y(\$genblock$spm.v:14$12[12].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _244_
  (
    .A1(_056_),
    .A2(_060_),
    .B1(_058_),
    .Y(_219_)
  );


  sky130_fd_sc_hd__inv_1
  _245_
  (
    .A(rst),
    .Y(_220_)
  );


  sky130_fd_sc_hd__inv_1
  _246_
  (
    .A(rst),
    .Y(_221_)
  );


  sky130_fd_sc_hd__nand2_1
  _247_
  (
    .A(y),
    .B(x[13]),
    .Y(_063_)
  );


  sky130_fd_sc_hd__nand2_1
  _248_
  (
    .A(\$genblock$spm.v:14$13[13].csa.sc ),
    .B(\$genblock$spm.v:14$14[14].csa.sum ),
    .Y(_064_)
  );


  sky130_fd_sc_hd__nor2_1
  _249_
  (
    .A(\$genblock$spm.v:14$13[13].csa.sc ),
    .B(\$genblock$spm.v:14$14[14].csa.sum ),
    .Y(_066_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _250_
  (
    .A(_064_),
    .SLEEP(_066_),
    .X(_068_)
  );


  sky130_fd_sc_hd__xnor2_1
  _251_
  (
    .A(_063_),
    .B(_068_),
    .Y(\$genblock$spm.v:14$13[13].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _252_
  (
    .A1(_063_),
    .A2(_066_),
    .B1(_064_),
    .Y(_222_)
  );


  sky130_fd_sc_hd__inv_1
  _253_
  (
    .A(rst),
    .Y(_001_)
  );


  sky130_fd_sc_hd__inv_1
  _254_
  (
    .A(rst),
    .Y(_002_)
  );


  sky130_fd_sc_hd__nand2_1
  _255_
  (
    .A(y),
    .B(x[14]),
    .Y(_070_)
  );


  sky130_fd_sc_hd__nand2_1
  _256_
  (
    .A(\$genblock$spm.v:14$14[14].csa.sc ),
    .B(\$genblock$spm.v:14$15[15].csa.sum ),
    .Y(_071_)
  );


  sky130_fd_sc_hd__nor2_1
  _257_
  (
    .A(\$genblock$spm.v:14$14[14].csa.sc ),
    .B(\$genblock$spm.v:14$15[15].csa.sum ),
    .Y(_072_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _258_
  (
    .A(_071_),
    .SLEEP(_072_),
    .X(_074_)
  );


  sky130_fd_sc_hd__xnor2_1
  _259_
  (
    .A(_070_),
    .B(_074_),
    .Y(\$genblock$spm.v:14$14[14].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _260_
  (
    .A1(_070_),
    .A2(_072_),
    .B1(_071_),
    .Y(_003_)
  );


  sky130_fd_sc_hd__inv_1
  _261_
  (
    .A(rst),
    .Y(_004_)
  );


  sky130_fd_sc_hd__inv_1
  _262_
  (
    .A(rst),
    .Y(_005_)
  );


  sky130_fd_sc_hd__nand2_1
  _263_
  (
    .A(y),
    .B(x[15]),
    .Y(_077_)
  );


  sky130_fd_sc_hd__nand2_1
  _264_
  (
    .A(\$genblock$spm.v:14$15[15].csa.sc ),
    .B(\$genblock$spm.v:14$16[16].csa.sum ),
    .Y(_078_)
  );


  sky130_fd_sc_hd__nor2_1
  _265_
  (
    .A(\$genblock$spm.v:14$15[15].csa.sc ),
    .B(\$genblock$spm.v:14$16[16].csa.sum ),
    .Y(_079_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _266_
  (
    .A(_078_),
    .SLEEP(_079_),
    .X(_080_)
  );


  sky130_fd_sc_hd__xnor2_1
  _267_
  (
    .A(_077_),
    .B(_080_),
    .Y(\$genblock$spm.v:14$15[15].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _268_
  (
    .A1(_077_),
    .A2(_079_),
    .B1(_078_),
    .Y(_006_)
  );


  sky130_fd_sc_hd__inv_1
  _269_
  (
    .A(rst),
    .Y(_007_)
  );


  sky130_fd_sc_hd__inv_1
  _270_
  (
    .A(rst),
    .Y(_008_)
  );


  sky130_fd_sc_hd__nand2_1
  _271_
  (
    .A(y),
    .B(x[16]),
    .Y(_084_)
  );


  sky130_fd_sc_hd__nand2_1
  _272_
  (
    .A(\$genblock$spm.v:14$16[16].csa.sc ),
    .B(\$genblock$spm.v:14$17[17].csa.sum ),
    .Y(_085_)
  );


  sky130_fd_sc_hd__nor2_1
  _273_
  (
    .A(\$genblock$spm.v:14$16[16].csa.sc ),
    .B(\$genblock$spm.v:14$17[17].csa.sum ),
    .Y(_086_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _274_
  (
    .A(_085_),
    .SLEEP(_086_),
    .X(_087_)
  );


  sky130_fd_sc_hd__xnor2_1
  _275_
  (
    .A(_084_),
    .B(_087_),
    .Y(\$genblock$spm.v:14$16[16].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _276_
  (
    .A1(_084_),
    .A2(_086_),
    .B1(_085_),
    .Y(_009_)
  );


  sky130_fd_sc_hd__inv_1
  _277_
  (
    .A(rst),
    .Y(_010_)
  );


  sky130_fd_sc_hd__inv_1
  _278_
  (
    .A(rst),
    .Y(_011_)
  );


  sky130_fd_sc_hd__nand2_1
  _279_
  (
    .A(y),
    .B(x[17]),
    .Y(_091_)
  );


  sky130_fd_sc_hd__nand2_1
  _280_
  (
    .A(\$genblock$spm.v:14$17[17].csa.sc ),
    .B(\$genblock$spm.v:14$18[18].csa.sum ),
    .Y(_092_)
  );


  sky130_fd_sc_hd__nor2_1
  _281_
  (
    .A(\$genblock$spm.v:14$17[17].csa.sc ),
    .B(\$genblock$spm.v:14$18[18].csa.sum ),
    .Y(_093_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _282_
  (
    .A(_092_),
    .SLEEP(_093_),
    .X(_094_)
  );


  sky130_fd_sc_hd__xnor2_1
  _283_
  (
    .A(_091_),
    .B(_094_),
    .Y(\$genblock$spm.v:14$17[17].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _284_
  (
    .A1(_091_),
    .A2(_093_),
    .B1(_092_),
    .Y(_012_)
  );


  sky130_fd_sc_hd__inv_1
  _285_
  (
    .A(rst),
    .Y(_013_)
  );


  sky130_fd_sc_hd__inv_1
  _286_
  (
    .A(rst),
    .Y(_014_)
  );


  sky130_fd_sc_hd__nand2_1
  _287_
  (
    .A(y),
    .B(x[18]),
    .Y(_098_)
  );


  sky130_fd_sc_hd__nand2_1
  _288_
  (
    .A(\$genblock$spm.v:14$18[18].csa.sc ),
    .B(\$genblock$spm.v:14$19[19].csa.sum ),
    .Y(_099_)
  );


  sky130_fd_sc_hd__nor2_1
  _289_
  (
    .A(\$genblock$spm.v:14$18[18].csa.sc ),
    .B(\$genblock$spm.v:14$19[19].csa.sum ),
    .Y(_100_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _290_
  (
    .A(_099_),
    .SLEEP(_100_),
    .X(_101_)
  );


  sky130_fd_sc_hd__xnor2_1
  _291_
  (
    .A(_098_),
    .B(_101_),
    .Y(\$genblock$spm.v:14$18[18].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _292_
  (
    .A1(_098_),
    .A2(_100_),
    .B1(_099_),
    .Y(_015_)
  );


  sky130_fd_sc_hd__inv_1
  _293_
  (
    .A(rst),
    .Y(_016_)
  );


  sky130_fd_sc_hd__inv_1
  _294_
  (
    .A(rst),
    .Y(_017_)
  );


  sky130_fd_sc_hd__nand2_1
  _295_
  (
    .A(y),
    .B(x[19]),
    .Y(_104_)
  );


  sky130_fd_sc_hd__nand2_1
  _296_
  (
    .A(\$genblock$spm.v:14$19[19].csa.sc ),
    .B(\$genblock$spm.v:14$20[20].csa.sum ),
    .Y(_106_)
  );


  sky130_fd_sc_hd__nor2_1
  _297_
  (
    .A(\$genblock$spm.v:14$19[19].csa.sc ),
    .B(\$genblock$spm.v:14$20[20].csa.sum ),
    .Y(_107_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _298_
  (
    .A(_106_),
    .SLEEP(_107_),
    .X(_108_)
  );


  sky130_fd_sc_hd__xnor2_1
  _299_
  (
    .A(_104_),
    .B(_108_),
    .Y(\$genblock$spm.v:14$19[19].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _300_
  (
    .A1(_104_),
    .A2(_107_),
    .B1(_106_),
    .Y(_018_)
  );


  sky130_fd_sc_hd__inv_1
  _301_
  (
    .A(rst),
    .Y(_019_)
  );


  sky130_fd_sc_hd__inv_1
  _302_
  (
    .A(rst),
    .Y(_020_)
  );


  sky130_fd_sc_hd__nand2_1
  _303_
  (
    .A(y),
    .B(x[1]),
    .Y(_110_)
  );


  sky130_fd_sc_hd__nand2_1
  _304_
  (
    .A(\$genblock$spm.v:14$1[1].csa.sc ),
    .B(\$genblock$spm.v:14$2[2].csa.sum ),
    .Y(_112_)
  );


  sky130_fd_sc_hd__nor2_1
  _305_
  (
    .A(\$genblock$spm.v:14$1[1].csa.sc ),
    .B(\$genblock$spm.v:14$2[2].csa.sum ),
    .Y(_114_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _306_
  (
    .A(_112_),
    .SLEEP(_114_),
    .X(_115_)
  );


  sky130_fd_sc_hd__xnor2_1
  _307_
  (
    .A(_110_),
    .B(_115_),
    .Y(\$genblock$spm.v:14$1[1].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _308_
  (
    .A1(_110_),
    .A2(_114_),
    .B1(_112_),
    .Y(_021_)
  );


  sky130_fd_sc_hd__inv_1
  _309_
  (
    .A(rst),
    .Y(_022_)
  );


  sky130_fd_sc_hd__inv_1
  _310_
  (
    .A(rst),
    .Y(_023_)
  );


  sky130_fd_sc_hd__nand2_1
  _311_
  (
    .A(y),
    .B(x[20]),
    .Y(_116_)
  );


  sky130_fd_sc_hd__nand2_1
  _312_
  (
    .A(\$genblock$spm.v:14$20[20].csa.sc ),
    .B(\$genblock$spm.v:14$21[21].csa.sum ),
    .Y(_118_)
  );


  sky130_fd_sc_hd__nor2_1
  _313_
  (
    .A(\$genblock$spm.v:14$20[20].csa.sc ),
    .B(\$genblock$spm.v:14$21[21].csa.sum ),
    .Y(_120_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _314_
  (
    .A(_118_),
    .SLEEP(_120_),
    .X(_122_)
  );


  sky130_fd_sc_hd__xnor2_1
  _315_
  (
    .A(_116_),
    .B(_122_),
    .Y(\$genblock$spm.v:14$20[20].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _316_
  (
    .A1(_116_),
    .A2(_120_),
    .B1(_118_),
    .Y(_024_)
  );


  sky130_fd_sc_hd__inv_1
  _317_
  (
    .A(rst),
    .Y(_025_)
  );


  sky130_fd_sc_hd__inv_1
  _318_
  (
    .A(rst),
    .Y(_026_)
  );


  sky130_fd_sc_hd__nand2_1
  _319_
  (
    .A(y),
    .B(x[21]),
    .Y(_123_)
  );


  sky130_fd_sc_hd__nand2_1
  _320_
  (
    .A(\$genblock$spm.v:14$21[21].csa.sc ),
    .B(\$genblock$spm.v:14$22[22].csa.sum ),
    .Y(_124_)
  );


  sky130_fd_sc_hd__nor2_1
  _321_
  (
    .A(\$genblock$spm.v:14$21[21].csa.sc ),
    .B(\$genblock$spm.v:14$22[22].csa.sum ),
    .Y(_126_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _322_
  (
    .A(_124_),
    .SLEEP(_126_),
    .X(_128_)
  );


  sky130_fd_sc_hd__xnor2_1
  _323_
  (
    .A(_123_),
    .B(_128_),
    .Y(\$genblock$spm.v:14$21[21].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _324_
  (
    .A1(_123_),
    .A2(_126_),
    .B1(_124_),
    .Y(_027_)
  );


  sky130_fd_sc_hd__inv_1
  _325_
  (
    .A(rst),
    .Y(_028_)
  );


  sky130_fd_sc_hd__inv_1
  _326_
  (
    .A(rst),
    .Y(_029_)
  );


  sky130_fd_sc_hd__nand2_1
  _327_
  (
    .A(y),
    .B(x[22]),
    .Y(_130_)
  );


  sky130_fd_sc_hd__nand2_1
  _328_
  (
    .A(\$genblock$spm.v:14$22[22].csa.sc ),
    .B(\$genblock$spm.v:14$23[23].csa.sum ),
    .Y(_131_)
  );


  sky130_fd_sc_hd__nor2_1
  _329_
  (
    .A(\$genblock$spm.v:14$22[22].csa.sc ),
    .B(\$genblock$spm.v:14$23[23].csa.sum ),
    .Y(_132_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _330_
  (
    .A(_131_),
    .SLEEP(_132_),
    .X(_134_)
  );


  sky130_fd_sc_hd__xnor2_1
  _331_
  (
    .A(_130_),
    .B(_134_),
    .Y(\$genblock$spm.v:14$22[22].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _332_
  (
    .A1(_130_),
    .A2(_132_),
    .B1(_131_),
    .Y(_030_)
  );


  sky130_fd_sc_hd__inv_1
  _333_
  (
    .A(rst),
    .Y(_031_)
  );


  sky130_fd_sc_hd__inv_1
  _334_
  (
    .A(rst),
    .Y(_032_)
  );


  sky130_fd_sc_hd__nand2_1
  _335_
  (
    .A(y),
    .B(x[23]),
    .Y(_137_)
  );


  sky130_fd_sc_hd__nand2_1
  _336_
  (
    .A(\$genblock$spm.v:14$23[23].csa.sc ),
    .B(\$genblock$spm.v:14$24[24].csa.sum ),
    .Y(_138_)
  );


  sky130_fd_sc_hd__nor2_1
  _337_
  (
    .A(\$genblock$spm.v:14$23[23].csa.sc ),
    .B(\$genblock$spm.v:14$24[24].csa.sum ),
    .Y(_139_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _338_
  (
    .A(_138_),
    .SLEEP(_139_),
    .X(_140_)
  );


  sky130_fd_sc_hd__xnor2_1
  _339_
  (
    .A(_137_),
    .B(_140_),
    .Y(\$genblock$spm.v:14$23[23].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _340_
  (
    .A1(_137_),
    .A2(_139_),
    .B1(_138_),
    .Y(_033_)
  );


  sky130_fd_sc_hd__inv_1
  _341_
  (
    .A(rst),
    .Y(_034_)
  );


  sky130_fd_sc_hd__inv_1
  _342_
  (
    .A(rst),
    .Y(_035_)
  );


  sky130_fd_sc_hd__nand2_1
  _343_
  (
    .A(y),
    .B(x[24]),
    .Y(_145_)
  );


  sky130_fd_sc_hd__nand2_1
  _344_
  (
    .A(\$genblock$spm.v:14$24[24].csa.sc ),
    .B(\$genblock$spm.v:14$25[25].csa.sum ),
    .Y(_147_)
  );


  sky130_fd_sc_hd__nor2_1
  _345_
  (
    .A(\$genblock$spm.v:14$24[24].csa.sc ),
    .B(\$genblock$spm.v:14$25[25].csa.sum ),
    .Y(_149_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _346_
  (
    .A(_147_),
    .SLEEP(_149_),
    .X(_151_)
  );


  sky130_fd_sc_hd__xnor2_1
  _347_
  (
    .A(_145_),
    .B(_151_),
    .Y(\$genblock$spm.v:14$24[24].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _348_
  (
    .A1(_145_),
    .A2(_149_),
    .B1(_147_),
    .Y(_036_)
  );


  sky130_fd_sc_hd__inv_1
  _349_
  (
    .A(rst),
    .Y(_037_)
  );


  sky130_fd_sc_hd__inv_1
  _350_
  (
    .A(rst),
    .Y(_038_)
  );


  sky130_fd_sc_hd__nand2_1
  _351_
  (
    .A(y),
    .B(x[25]),
    .Y(_152_)
  );


  sky130_fd_sc_hd__nand2_1
  _352_
  (
    .A(\$genblock$spm.v:14$25[25].csa.sc ),
    .B(\$genblock$spm.v:14$26[26].csa.sum ),
    .Y(_153_)
  );


  sky130_fd_sc_hd__nor2_1
  _353_
  (
    .A(\$genblock$spm.v:14$25[25].csa.sc ),
    .B(\$genblock$spm.v:14$26[26].csa.sum ),
    .Y(_154_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _354_
  (
    .A(_153_),
    .SLEEP(_154_),
    .X(_155_)
  );


  sky130_fd_sc_hd__xnor2_1
  _355_
  (
    .A(_152_),
    .B(_155_),
    .Y(\$genblock$spm.v:14$25[25].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _356_
  (
    .A1(_152_),
    .A2(_154_),
    .B1(_153_),
    .Y(_039_)
  );


  sky130_fd_sc_hd__inv_1
  _357_
  (
    .A(rst),
    .Y(_040_)
  );


  sky130_fd_sc_hd__inv_1
  _358_
  (
    .A(rst),
    .Y(_041_)
  );


  sky130_fd_sc_hd__nand2_1
  _359_
  (
    .A(y),
    .B(x[26]),
    .Y(_156_)
  );


  sky130_fd_sc_hd__nand2_1
  _360_
  (
    .A(\$genblock$spm.v:14$26[26].csa.sc ),
    .B(\$genblock$spm.v:14$27[27].csa.sum ),
    .Y(_157_)
  );


  sky130_fd_sc_hd__nor2_1
  _361_
  (
    .A(\$genblock$spm.v:14$26[26].csa.sc ),
    .B(\$genblock$spm.v:14$27[27].csa.sum ),
    .Y(_158_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _362_
  (
    .A(_157_),
    .SLEEP(_158_),
    .X(_159_)
  );


  sky130_fd_sc_hd__xnor2_1
  _363_
  (
    .A(_156_),
    .B(_159_),
    .Y(\$genblock$spm.v:14$26[26].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _364_
  (
    .A1(_156_),
    .A2(_158_),
    .B1(_157_),
    .Y(_042_)
  );


  sky130_fd_sc_hd__inv_1
  _365_
  (
    .A(rst),
    .Y(_043_)
  );


  sky130_fd_sc_hd__inv_1
  _366_
  (
    .A(rst),
    .Y(_044_)
  );


  sky130_fd_sc_hd__nand2_1
  _367_
  (
    .A(y),
    .B(x[27]),
    .Y(_160_)
  );


  sky130_fd_sc_hd__nand2_1
  _368_
  (
    .A(\$genblock$spm.v:14$27[27].csa.sc ),
    .B(\$genblock$spm.v:14$28[28].csa.sum ),
    .Y(_161_)
  );


  sky130_fd_sc_hd__nor2_1
  _369_
  (
    .A(\$genblock$spm.v:14$27[27].csa.sc ),
    .B(\$genblock$spm.v:14$28[28].csa.sum ),
    .Y(_162_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _370_
  (
    .A(_161_),
    .SLEEP(_162_),
    .X(_163_)
  );


  sky130_fd_sc_hd__xnor2_1
  _371_
  (
    .A(_160_),
    .B(_163_),
    .Y(\$genblock$spm.v:14$27[27].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _372_
  (
    .A1(_160_),
    .A2(_162_),
    .B1(_161_),
    .Y(_049_)
  );


  sky130_fd_sc_hd__inv_1
  _373_
  (
    .A(rst),
    .Y(_051_)
  );


  sky130_fd_sc_hd__inv_1
  _374_
  (
    .A(rst),
    .Y(_053_)
  );


  sky130_fd_sc_hd__nand2_1
  _375_
  (
    .A(y),
    .B(x[28]),
    .Y(_164_)
  );


  sky130_fd_sc_hd__nand2_1
  _376_
  (
    .A(\$genblock$spm.v:14$28[28].csa.sc ),
    .B(\$genblock$spm.v:14$29[29].csa.sum ),
    .Y(_165_)
  );


  sky130_fd_sc_hd__nor2_1
  _377_
  (
    .A(\$genblock$spm.v:14$28[28].csa.sc ),
    .B(\$genblock$spm.v:14$29[29].csa.sum ),
    .Y(_166_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _378_
  (
    .A(_165_),
    .SLEEP(_166_),
    .X(_167_)
  );


  sky130_fd_sc_hd__xnor2_1
  _379_
  (
    .A(_164_),
    .B(_167_),
    .Y(\$genblock$spm.v:14$28[28].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _380_
  (
    .A1(_164_),
    .A2(_166_),
    .B1(_165_),
    .Y(_057_)
  );


  sky130_fd_sc_hd__inv_1
  _381_
  (
    .A(rst),
    .Y(_059_)
  );


  sky130_fd_sc_hd__inv_1
  _382_
  (
    .A(rst),
    .Y(_061_)
  );


  sky130_fd_sc_hd__nand2_1
  _383_
  (
    .A(y),
    .B(x[29]),
    .Y(_168_)
  );


  sky130_fd_sc_hd__nand2_1
  _384_
  (
    .A(\$genblock$spm.v:14$29[29].csa.sc ),
    .B(\$genblock$spm.v:14$30[30].csa.sum ),
    .Y(_169_)
  );


  sky130_fd_sc_hd__nor2_1
  _385_
  (
    .A(\$genblock$spm.v:14$29[29].csa.sc ),
    .B(\$genblock$spm.v:14$30[30].csa.sum ),
    .Y(_170_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _386_
  (
    .A(_169_),
    .SLEEP(_170_),
    .X(_171_)
  );


  sky130_fd_sc_hd__xnor2_1
  _387_
  (
    .A(_168_),
    .B(_171_),
    .Y(\$genblock$spm.v:14$29[29].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _388_
  (
    .A1(_168_),
    .A2(_170_),
    .B1(_169_),
    .Y(_065_)
  );


  sky130_fd_sc_hd__inv_1
  _389_
  (
    .A(rst),
    .Y(_067_)
  );


  sky130_fd_sc_hd__inv_1
  _390_
  (
    .A(rst),
    .Y(_069_)
  );


  sky130_fd_sc_hd__nand2_1
  _391_
  (
    .A(y),
    .B(x[2]),
    .Y(_172_)
  );


  sky130_fd_sc_hd__nand2_1
  _392_
  (
    .A(\$genblock$spm.v:14$2[2].csa.sc ),
    .B(\$genblock$spm.v:14$3[3].csa.sum ),
    .Y(_173_)
  );


  sky130_fd_sc_hd__nor2_1
  _393_
  (
    .A(\$genblock$spm.v:14$2[2].csa.sc ),
    .B(\$genblock$spm.v:14$3[3].csa.sum ),
    .Y(_174_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _394_
  (
    .A(_173_),
    .SLEEP(_174_),
    .X(_175_)
  );


  sky130_fd_sc_hd__xnor2_1
  _395_
  (
    .A(_172_),
    .B(_175_),
    .Y(\$genblock$spm.v:14$2[2].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _396_
  (
    .A1(_172_),
    .A2(_174_),
    .B1(_173_),
    .Y(_073_)
  );


  sky130_fd_sc_hd__inv_1
  _397_
  (
    .A(rst),
    .Y(_075_)
  );


  sky130_fd_sc_hd__inv_1
  _398_
  (
    .A(rst),
    .Y(_076_)
  );


  sky130_fd_sc_hd__nand2_1
  _399_
  (
    .A(y),
    .B(x[30]),
    .Y(_176_)
  );


  sky130_fd_sc_hd__nand2_1
  _400_
  (
    .A(\$genblock$spm.v:14$30[30].csa.sc ),
    .B(\tcmp.s ),
    .Y(_177_)
  );


  sky130_fd_sc_hd__nor2_1
  _401_
  (
    .A(\$genblock$spm.v:14$30[30].csa.sc ),
    .B(\tcmp.s ),
    .Y(_178_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _402_
  (
    .A(_177_),
    .SLEEP(_178_),
    .X(_179_)
  );


  sky130_fd_sc_hd__xnor2_1
  _403_
  (
    .A(_176_),
    .B(_179_),
    .Y(\$genblock$spm.v:14$30[30].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _404_
  (
    .A1(_176_),
    .A2(_178_),
    .B1(_177_),
    .Y(_081_)
  );


  sky130_fd_sc_hd__inv_1
  _405_
  (
    .A(rst),
    .Y(_082_)
  );


  sky130_fd_sc_hd__inv_1
  _406_
  (
    .A(rst),
    .Y(_083_)
  );


  sky130_fd_sc_hd__nand2_1
  _407_
  (
    .A(y),
    .B(x[3]),
    .Y(_180_)
  );


  sky130_fd_sc_hd__nand2_1
  _408_
  (
    .A(\$genblock$spm.v:14$3[3].csa.sc ),
    .B(\$genblock$spm.v:14$4[4].csa.sum ),
    .Y(_181_)
  );


  sky130_fd_sc_hd__nor2_1
  _409_
  (
    .A(\$genblock$spm.v:14$3[3].csa.sc ),
    .B(\$genblock$spm.v:14$4[4].csa.sum ),
    .Y(_182_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _410_
  (
    .A(_181_),
    .SLEEP(_182_),
    .X(_183_)
  );


  sky130_fd_sc_hd__xnor2_1
  _411_
  (
    .A(_180_),
    .B(_183_),
    .Y(\$genblock$spm.v:14$3[3].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _412_
  (
    .A1(_180_),
    .A2(_182_),
    .B1(_181_),
    .Y(_088_)
  );


  sky130_fd_sc_hd__inv_1
  _413_
  (
    .A(rst),
    .Y(_089_)
  );


  sky130_fd_sc_hd__inv_1
  _414_
  (
    .A(rst),
    .Y(_090_)
  );


  sky130_fd_sc_hd__nand2_1
  _415_
  (
    .A(y),
    .B(x[4]),
    .Y(_184_)
  );


  sky130_fd_sc_hd__nand2_1
  _416_
  (
    .A(\$genblock$spm.v:14$4[4].csa.sc ),
    .B(\$genblock$spm.v:14$5[5].csa.sum ),
    .Y(_185_)
  );


  sky130_fd_sc_hd__nor2_1
  _417_
  (
    .A(\$genblock$spm.v:14$4[4].csa.sc ),
    .B(\$genblock$spm.v:14$5[5].csa.sum ),
    .Y(_186_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _418_
  (
    .A(_185_),
    .SLEEP(_186_),
    .X(_187_)
  );


  sky130_fd_sc_hd__xnor2_1
  _419_
  (
    .A(_184_),
    .B(_187_),
    .Y(\$genblock$spm.v:14$4[4].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _420_
  (
    .A1(_184_),
    .A2(_186_),
    .B1(_185_),
    .Y(_095_)
  );


  sky130_fd_sc_hd__inv_1
  _421_
  (
    .A(rst),
    .Y(_096_)
  );


  sky130_fd_sc_hd__inv_1
  _422_
  (
    .A(rst),
    .Y(_097_)
  );


  sky130_fd_sc_hd__nand2_1
  _423_
  (
    .A(y),
    .B(x[5]),
    .Y(_188_)
  );


  sky130_fd_sc_hd__nand2_1
  _424_
  (
    .A(\$genblock$spm.v:14$5[5].csa.sc ),
    .B(\$genblock$spm.v:14$6[6].csa.sum ),
    .Y(_189_)
  );


  sky130_fd_sc_hd__nor2_1
  _425_
  (
    .A(\$genblock$spm.v:14$5[5].csa.sc ),
    .B(\$genblock$spm.v:14$6[6].csa.sum ),
    .Y(_190_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _426_
  (
    .A(_189_),
    .SLEEP(_190_),
    .X(_191_)
  );


  sky130_fd_sc_hd__xnor2_1
  _427_
  (
    .A(_188_),
    .B(_191_),
    .Y(\$genblock$spm.v:14$5[5].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _428_
  (
    .A1(_188_),
    .A2(_190_),
    .B1(_189_),
    .Y(_102_)
  );


  sky130_fd_sc_hd__inv_1
  _429_
  (
    .A(rst),
    .Y(_103_)
  );


  sky130_fd_sc_hd__inv_1
  _430_
  (
    .A(rst),
    .Y(_105_)
  );


  sky130_fd_sc_hd__nand2_1
  _431_
  (
    .A(y),
    .B(x[6]),
    .Y(_192_)
  );


  sky130_fd_sc_hd__nand2_1
  _432_
  (
    .A(\$genblock$spm.v:14$6[6].csa.sc ),
    .B(\$genblock$spm.v:14$7[7].csa.sum ),
    .Y(_193_)
  );


  sky130_fd_sc_hd__nor2_1
  _433_
  (
    .A(\$genblock$spm.v:14$6[6].csa.sc ),
    .B(\$genblock$spm.v:14$7[7].csa.sum ),
    .Y(_194_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _434_
  (
    .A(_193_),
    .SLEEP(_194_),
    .X(_195_)
  );


  sky130_fd_sc_hd__xnor2_1
  _435_
  (
    .A(_192_),
    .B(_195_),
    .Y(\$genblock$spm.v:14$6[6].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _436_
  (
    .A1(_192_),
    .A2(_194_),
    .B1(_193_),
    .Y(_109_)
  );


  sky130_fd_sc_hd__inv_1
  _437_
  (
    .A(rst),
    .Y(_111_)
  );


  sky130_fd_sc_hd__inv_1
  _438_
  (
    .A(rst),
    .Y(_113_)
  );


  sky130_fd_sc_hd__nand2_1
  _439_
  (
    .A(y),
    .B(x[7]),
    .Y(_196_)
  );


  sky130_fd_sc_hd__nand2_1
  _440_
  (
    .A(\$genblock$spm.v:14$7[7].csa.sc ),
    .B(\$genblock$spm.v:14$8[8].csa.sum ),
    .Y(_197_)
  );


  sky130_fd_sc_hd__nor2_1
  _441_
  (
    .A(\$genblock$spm.v:14$7[7].csa.sc ),
    .B(\$genblock$spm.v:14$8[8].csa.sum ),
    .Y(_198_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _442_
  (
    .A(_197_),
    .SLEEP(_198_),
    .X(_199_)
  );


  sky130_fd_sc_hd__xnor2_1
  _443_
  (
    .A(_196_),
    .B(_199_),
    .Y(\$genblock$spm.v:14$7[7].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _444_
  (
    .A1(_196_),
    .A2(_198_),
    .B1(_197_),
    .Y(_117_)
  );


  sky130_fd_sc_hd__inv_1
  _445_
  (
    .A(rst),
    .Y(_119_)
  );


  sky130_fd_sc_hd__inv_1
  _446_
  (
    .A(rst),
    .Y(_121_)
  );


  sky130_fd_sc_hd__nand2_1
  _447_
  (
    .A(y),
    .B(x[8]),
    .Y(_200_)
  );


  sky130_fd_sc_hd__nand2_1
  _448_
  (
    .A(\$genblock$spm.v:14$8[8].csa.sc ),
    .B(\$genblock$spm.v:14$9[9].csa.sum ),
    .Y(_201_)
  );


  sky130_fd_sc_hd__nor2_1
  _449_
  (
    .A(\$genblock$spm.v:14$8[8].csa.sc ),
    .B(\$genblock$spm.v:14$9[9].csa.sum ),
    .Y(_202_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _450_
  (
    .A(_201_),
    .SLEEP(_202_),
    .X(_203_)
  );


  sky130_fd_sc_hd__xnor2_1
  _451_
  (
    .A(_200_),
    .B(_203_),
    .Y(\$genblock$spm.v:14$8[8].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _452_
  (
    .A1(_200_),
    .A2(_202_),
    .B1(_201_),
    .Y(_125_)
  );


  sky130_fd_sc_hd__inv_1
  _453_
  (
    .A(rst),
    .Y(_127_)
  );


  sky130_fd_sc_hd__inv_1
  _454_
  (
    .A(rst),
    .Y(_129_)
  );


  sky130_fd_sc_hd__nand2_1
  _455_
  (
    .A(y),
    .B(x[9]),
    .Y(_204_)
  );


  sky130_fd_sc_hd__nand2_1
  _456_
  (
    .A(\$genblock$spm.v:14$9[9].csa.sc ),
    .B(\$genblock$spm.v:14$10[10].csa.sum ),
    .Y(_205_)
  );


  sky130_fd_sc_hd__nor2_1
  _457_
  (
    .A(\$genblock$spm.v:14$9[9].csa.sc ),
    .B(\$genblock$spm.v:14$10[10].csa.sum ),
    .Y(_206_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _458_
  (
    .A(_205_),
    .SLEEP(_206_),
    .X(_207_)
  );


  sky130_fd_sc_hd__xnor2_1
  _459_
  (
    .A(_204_),
    .B(_207_),
    .Y(\$genblock$spm.v:14$9[9].csa.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _460_
  (
    .A1(_204_),
    .A2(_206_),
    .B1(_205_),
    .Y(_133_)
  );


  sky130_fd_sc_hd__inv_1
  _461_
  (
    .A(rst),
    .Y(_135_)
  );


  sky130_fd_sc_hd__inv_1
  _462_
  (
    .A(rst),
    .Y(_136_)
  );


  sky130_fd_sc_hd__nand2_1
  _463_
  (
    .A(y),
    .B(x[0]),
    .Y(_208_)
  );


  sky130_fd_sc_hd__nand2_1
  _464_
  (
    .A(\csa0.sc ),
    .B(\$genblock$spm.v:14$1[1].csa.sum ),
    .Y(_209_)
  );


  sky130_fd_sc_hd__nor2_1
  _465_
  (
    .A(\csa0.sc ),
    .B(\$genblock$spm.v:14$1[1].csa.sum ),
    .Y(_210_)
  );


  sky130_fd_sc_hd__lpflow_isobufsrc_1
  _466_
  (
    .A(_209_),
    .SLEEP(_210_),
    .X(_211_)
  );


  sky130_fd_sc_hd__xnor2_1
  _467_
  (
    .A(_208_),
    .B(_211_),
    .Y(\csa0.hsum2 )
  );


  sky130_fd_sc_hd__o21ai_0
  _468_
  (
    .A1(_208_),
    .A2(_210_),
    .B1(_209_),
    .Y(_141_)
  );


  sky130_fd_sc_hd__inv_1
  _469_
  (
    .A(rst),
    .Y(_142_)
  );


  sky130_fd_sc_hd__inv_1
  _470_
  (
    .A(rst),
    .Y(_143_)
  );


  sky130_fd_sc_hd__nand2_1
  _471_
  (
    .A(x[31]),
    .B(y),
    .Y(_212_)
  );


  sky130_fd_sc_hd__inv_1
  _472_
  (
    .A(\tcmp.z ),
    .Y(_213_)
  );


  sky130_fd_sc_hd__nand2_1
  _473_
  (
    .A(_212_),
    .B(_213_),
    .Y(_144_)
  );


  sky130_fd_sc_hd__xnor2_1
  _474_
  (
    .A(\tcmp.z ),
    .B(_212_),
    .Y(_146_)
  );


  sky130_fd_sc_hd__inv_1
  _475_
  (
    .A(rst),
    .Y(_148_)
  );


  sky130_fd_sc_hd__inv_1
  _476_
  (
    .A(rst),
    .Y(_150_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _477_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$10[10].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$10[10].csa.sum ),
    .RESET_B(_215_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _478_
  (
    .CLK(clk),
    .D(_214_),
    .Q(\$genblock$spm.v:14$10[10].csa.sc ),
    .RESET_B(_217_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _479_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$11[11].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$11[11].csa.sum ),
    .RESET_B(_218_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _480_
  (
    .CLK(clk),
    .D(_216_),
    .Q(\$genblock$spm.v:14$11[11].csa.sc ),
    .RESET_B(_220_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _481_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$12[12].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$12[12].csa.sum ),
    .RESET_B(_221_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _482_
  (
    .CLK(clk),
    .D(_219_),
    .Q(\$genblock$spm.v:14$12[12].csa.sc ),
    .RESET_B(_001_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _483_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$13[13].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$13[13].csa.sum ),
    .RESET_B(_002_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _484_
  (
    .CLK(clk),
    .D(_222_),
    .Q(\$genblock$spm.v:14$13[13].csa.sc ),
    .RESET_B(_004_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _485_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$14[14].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$14[14].csa.sum ),
    .RESET_B(_005_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _486_
  (
    .CLK(clk),
    .D(_003_),
    .Q(\$genblock$spm.v:14$14[14].csa.sc ),
    .RESET_B(_007_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _487_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$15[15].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$15[15].csa.sum ),
    .RESET_B(_008_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _488_
  (
    .CLK(clk),
    .D(_006_),
    .Q(\$genblock$spm.v:14$15[15].csa.sc ),
    .RESET_B(_010_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _489_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$16[16].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$16[16].csa.sum ),
    .RESET_B(_011_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _490_
  (
    .CLK(clk),
    .D(_009_),
    .Q(\$genblock$spm.v:14$16[16].csa.sc ),
    .RESET_B(_013_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _491_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$17[17].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$17[17].csa.sum ),
    .RESET_B(_014_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _492_
  (
    .CLK(clk),
    .D(_012_),
    .Q(\$genblock$spm.v:14$17[17].csa.sc ),
    .RESET_B(_016_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _493_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$18[18].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$18[18].csa.sum ),
    .RESET_B(_017_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _494_
  (
    .CLK(clk),
    .D(_015_),
    .Q(\$genblock$spm.v:14$18[18].csa.sc ),
    .RESET_B(_019_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _495_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$19[19].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$19[19].csa.sum ),
    .RESET_B(_020_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _496_
  (
    .CLK(clk),
    .D(_018_),
    .Q(\$genblock$spm.v:14$19[19].csa.sc ),
    .RESET_B(_022_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _497_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$1[1].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$1[1].csa.sum ),
    .RESET_B(_023_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _498_
  (
    .CLK(clk),
    .D(_021_),
    .Q(\$genblock$spm.v:14$1[1].csa.sc ),
    .RESET_B(_025_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _499_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$20[20].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$20[20].csa.sum ),
    .RESET_B(_026_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _500_
  (
    .CLK(clk),
    .D(_024_),
    .Q(\$genblock$spm.v:14$20[20].csa.sc ),
    .RESET_B(_028_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _501_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$21[21].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$21[21].csa.sum ),
    .RESET_B(_029_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _502_
  (
    .CLK(clk),
    .D(_027_),
    .Q(\$genblock$spm.v:14$21[21].csa.sc ),
    .RESET_B(_031_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _503_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$22[22].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$22[22].csa.sum ),
    .RESET_B(_032_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _504_
  (
    .CLK(clk),
    .D(_030_),
    .Q(\$genblock$spm.v:14$22[22].csa.sc ),
    .RESET_B(_034_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _505_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$23[23].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$23[23].csa.sum ),
    .RESET_B(_035_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _506_
  (
    .CLK(clk),
    .D(_033_),
    .Q(\$genblock$spm.v:14$23[23].csa.sc ),
    .RESET_B(_037_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _507_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$24[24].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$24[24].csa.sum ),
    .RESET_B(_038_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _508_
  (
    .CLK(clk),
    .D(_036_),
    .Q(\$genblock$spm.v:14$24[24].csa.sc ),
    .RESET_B(_040_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _509_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$25[25].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$25[25].csa.sum ),
    .RESET_B(_041_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _510_
  (
    .CLK(clk),
    .D(_039_),
    .Q(\$genblock$spm.v:14$25[25].csa.sc ),
    .RESET_B(_043_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _511_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$26[26].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$26[26].csa.sum ),
    .RESET_B(_044_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _512_
  (
    .CLK(clk),
    .D(_042_),
    .Q(\$genblock$spm.v:14$26[26].csa.sc ),
    .RESET_B(_051_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _513_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$27[27].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$27[27].csa.sum ),
    .RESET_B(_053_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _514_
  (
    .CLK(clk),
    .D(_049_),
    .Q(\$genblock$spm.v:14$27[27].csa.sc ),
    .RESET_B(_059_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _515_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$28[28].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$28[28].csa.sum ),
    .RESET_B(_061_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _516_
  (
    .CLK(clk),
    .D(_057_),
    .Q(\$genblock$spm.v:14$28[28].csa.sc ),
    .RESET_B(_067_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _517_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$29[29].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$29[29].csa.sum ),
    .RESET_B(_069_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _518_
  (
    .CLK(clk),
    .D(_065_),
    .Q(\$genblock$spm.v:14$29[29].csa.sc ),
    .RESET_B(_075_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _519_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$2[2].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$2[2].csa.sum ),
    .RESET_B(_076_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _520_
  (
    .CLK(clk),
    .D(_073_),
    .Q(\$genblock$spm.v:14$2[2].csa.sc ),
    .RESET_B(_082_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _521_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$30[30].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$30[30].csa.sum ),
    .RESET_B(_083_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _522_
  (
    .CLK(clk),
    .D(_081_),
    .Q(\$genblock$spm.v:14$30[30].csa.sc ),
    .RESET_B(_089_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _523_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$3[3].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$3[3].csa.sum ),
    .RESET_B(_090_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _524_
  (
    .CLK(clk),
    .D(_088_),
    .Q(\$genblock$spm.v:14$3[3].csa.sc ),
    .RESET_B(_096_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _525_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$4[4].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$4[4].csa.sum ),
    .RESET_B(_097_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _526_
  (
    .CLK(clk),
    .D(_095_),
    .Q(\$genblock$spm.v:14$4[4].csa.sc ),
    .RESET_B(_103_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _527_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$5[5].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$5[5].csa.sum ),
    .RESET_B(_105_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _528_
  (
    .CLK(clk),
    .D(_102_),
    .Q(\$genblock$spm.v:14$5[5].csa.sc ),
    .RESET_B(_111_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _529_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$6[6].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$6[6].csa.sum ),
    .RESET_B(_113_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _530_
  (
    .CLK(clk),
    .D(_109_),
    .Q(\$genblock$spm.v:14$6[6].csa.sc ),
    .RESET_B(_119_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _531_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$7[7].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$7[7].csa.sum ),
    .RESET_B(_121_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _532_
  (
    .CLK(clk),
    .D(_117_),
    .Q(\$genblock$spm.v:14$7[7].csa.sc ),
    .RESET_B(_127_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _533_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$8[8].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$8[8].csa.sum ),
    .RESET_B(_129_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _534_
  (
    .CLK(clk),
    .D(_125_),
    .Q(\$genblock$spm.v:14$8[8].csa.sc ),
    .RESET_B(_135_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _535_
  (
    .CLK(clk),
    .D(\$genblock$spm.v:14$9[9].csa.hsum2 ),
    .Q(\$genblock$spm.v:14$9[9].csa.sum ),
    .RESET_B(_136_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _536_
  (
    .CLK(clk),
    .D(_133_),
    .Q(\$genblock$spm.v:14$9[9].csa.sc ),
    .RESET_B(_142_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _537_
  (
    .CLK(clk),
    .D(\csa0.hsum2 ),
    .Q(\csa0.sum ),
    .RESET_B(_143_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _538_
  (
    .CLK(clk),
    .D(_141_),
    .Q(\csa0.sc ),
    .RESET_B(_148_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _539_
  (
    .CLK(clk),
    .D(_146_),
    .Q(\tcmp.s ),
    .RESET_B(_150_)
  );


  sky130_fd_sc_hd__dfrtp_1
  _540_
  (
    .CLK(clk),
    .D(_144_),
    .Q(\tcmp.z ),
    .RESET_B(_000_)
  );

  assign \$genblock$spm.v:14$10[10].csa.clk  = clk;
  assign \$genblock$spm.v:14$10[10].csa.rst  = rst;
  assign \$genblock$spm.v:14$10[10].csa.y  = \$genblock$spm.v:14$11[11].csa.sum ;
  assign \$genblock$spm.v:14$11[11].csa.clk  = clk;
  assign \$genblock$spm.v:14$11[11].csa.rst  = rst;
  assign \$genblock$spm.v:14$11[11].csa.y  = \$genblock$spm.v:14$12[12].csa.sum ;
  assign \$genblock$spm.v:14$12[12].csa.clk  = clk;
  assign \$genblock$spm.v:14$12[12].csa.rst  = rst;
  assign \$genblock$spm.v:14$12[12].csa.y  = \$genblock$spm.v:14$13[13].csa.sum ;
  assign \$genblock$spm.v:14$13[13].csa.clk  = clk;
  assign \$genblock$spm.v:14$13[13].csa.rst  = rst;
  assign \$genblock$spm.v:14$13[13].csa.y  = \$genblock$spm.v:14$14[14].csa.sum ;
  assign \$genblock$spm.v:14$14[14].csa.clk  = clk;
  assign \$genblock$spm.v:14$14[14].csa.rst  = rst;
  assign \$genblock$spm.v:14$14[14].csa.y  = \$genblock$spm.v:14$15[15].csa.sum ;
  assign \$genblock$spm.v:14$15[15].csa.clk  = clk;
  assign \$genblock$spm.v:14$15[15].csa.rst  = rst;
  assign \$genblock$spm.v:14$15[15].csa.y  = \$genblock$spm.v:14$16[16].csa.sum ;
  assign \$genblock$spm.v:14$16[16].csa.clk  = clk;
  assign \$genblock$spm.v:14$16[16].csa.rst  = rst;
  assign \$genblock$spm.v:14$16[16].csa.y  = \$genblock$spm.v:14$17[17].csa.sum ;
  assign \$genblock$spm.v:14$17[17].csa.clk  = clk;
  assign \$genblock$spm.v:14$17[17].csa.rst  = rst;
  assign \$genblock$spm.v:14$17[17].csa.y  = \$genblock$spm.v:14$18[18].csa.sum ;
  assign \$genblock$spm.v:14$18[18].csa.clk  = clk;
  assign \$genblock$spm.v:14$18[18].csa.rst  = rst;
  assign \$genblock$spm.v:14$18[18].csa.y  = \$genblock$spm.v:14$19[19].csa.sum ;
  assign \$genblock$spm.v:14$19[19].csa.clk  = clk;
  assign \$genblock$spm.v:14$19[19].csa.rst  = rst;
  assign \$genblock$spm.v:14$19[19].csa.y  = \$genblock$spm.v:14$20[20].csa.sum ;
  assign \$genblock$spm.v:14$1[1].csa.clk  = clk;
  assign \$genblock$spm.v:14$1[1].csa.rst  = rst;
  assign \$genblock$spm.v:14$1[1].csa.y  = \$genblock$spm.v:14$2[2].csa.sum ;
  assign \$genblock$spm.v:14$20[20].csa.clk  = clk;
  assign \$genblock$spm.v:14$20[20].csa.rst  = rst;
  assign \$genblock$spm.v:14$20[20].csa.y  = \$genblock$spm.v:14$21[21].csa.sum ;
  assign \$genblock$spm.v:14$21[21].csa.clk  = clk;
  assign \$genblock$spm.v:14$21[21].csa.rst  = rst;
  assign \$genblock$spm.v:14$21[21].csa.y  = \$genblock$spm.v:14$22[22].csa.sum ;
  assign \$genblock$spm.v:14$22[22].csa.clk  = clk;
  assign \$genblock$spm.v:14$22[22].csa.rst  = rst;
  assign \$genblock$spm.v:14$22[22].csa.y  = \$genblock$spm.v:14$23[23].csa.sum ;
  assign \$genblock$spm.v:14$23[23].csa.clk  = clk;
  assign \$genblock$spm.v:14$23[23].csa.rst  = rst;
  assign \$genblock$spm.v:14$23[23].csa.y  = \$genblock$spm.v:14$24[24].csa.sum ;
  assign \$genblock$spm.v:14$24[24].csa.clk  = clk;
  assign \$genblock$spm.v:14$24[24].csa.rst  = rst;
  assign \$genblock$spm.v:14$24[24].csa.y  = \$genblock$spm.v:14$25[25].csa.sum ;
  assign \$genblock$spm.v:14$25[25].csa.clk  = clk;
  assign \$genblock$spm.v:14$25[25].csa.rst  = rst;
  assign \$genblock$spm.v:14$25[25].csa.y  = \$genblock$spm.v:14$26[26].csa.sum ;
  assign \$genblock$spm.v:14$26[26].csa.clk  = clk;
  assign \$genblock$spm.v:14$26[26].csa.rst  = rst;
  assign \$genblock$spm.v:14$26[26].csa.y  = \$genblock$spm.v:14$27[27].csa.sum ;
  assign \$genblock$spm.v:14$27[27].csa.clk  = clk;
  assign \$genblock$spm.v:14$27[27].csa.rst  = rst;
  assign \$genblock$spm.v:14$27[27].csa.y  = \$genblock$spm.v:14$28[28].csa.sum ;
  assign \$genblock$spm.v:14$28[28].csa.clk  = clk;
  assign \$genblock$spm.v:14$28[28].csa.rst  = rst;
  assign \$genblock$spm.v:14$28[28].csa.y  = \$genblock$spm.v:14$29[29].csa.sum ;
  assign \$genblock$spm.v:14$29[29].csa.clk  = clk;
  assign \$genblock$spm.v:14$29[29].csa.rst  = rst;
  assign \$genblock$spm.v:14$29[29].csa.y  = \$genblock$spm.v:14$30[30].csa.sum ;
  assign \$genblock$spm.v:14$2[2].csa.clk  = clk;
  assign \$genblock$spm.v:14$2[2].csa.rst  = rst;
  assign \$genblock$spm.v:14$2[2].csa.y  = \$genblock$spm.v:14$3[3].csa.sum ;
  assign \$genblock$spm.v:14$30[30].csa.clk  = clk;
  assign \$genblock$spm.v:14$30[30].csa.rst  = rst;
  assign \$genblock$spm.v:14$30[30].csa.y  = \tcmp.s ;
  assign \$genblock$spm.v:14$3[3].csa.clk  = clk;
  assign \$genblock$spm.v:14$3[3].csa.rst  = rst;
  assign \$genblock$spm.v:14$3[3].csa.y  = \$genblock$spm.v:14$4[4].csa.sum ;
  assign \$genblock$spm.v:14$4[4].csa.clk  = clk;
  assign \$genblock$spm.v:14$4[4].csa.rst  = rst;
  assign \$genblock$spm.v:14$4[4].csa.y  = \$genblock$spm.v:14$5[5].csa.sum ;
  assign \$genblock$spm.v:14$5[5].csa.clk  = clk;
  assign \$genblock$spm.v:14$5[5].csa.rst  = rst;
  assign \$genblock$spm.v:14$5[5].csa.y  = \$genblock$spm.v:14$6[6].csa.sum ;
  assign \$genblock$spm.v:14$6[6].csa.clk  = clk;
  assign \$genblock$spm.v:14$6[6].csa.rst  = rst;
  assign \$genblock$spm.v:14$6[6].csa.y  = \$genblock$spm.v:14$7[7].csa.sum ;
  assign \$genblock$spm.v:14$7[7].csa.clk  = clk;
  assign \$genblock$spm.v:14$7[7].csa.rst  = rst;
  assign \$genblock$spm.v:14$7[7].csa.y  = \$genblock$spm.v:14$8[8].csa.sum ;
  assign \$genblock$spm.v:14$8[8].csa.clk  = clk;
  assign \$genblock$spm.v:14$8[8].csa.rst  = rst;
  assign \$genblock$spm.v:14$8[8].csa.y  = \$genblock$spm.v:14$9[9].csa.sum ;
  assign \$genblock$spm.v:14$9[9].csa.clk  = clk;
  assign \$genblock$spm.v:14$9[9].csa.rst  = rst;
  assign \$genblock$spm.v:14$9[9].csa.y  = \$genblock$spm.v:14$10[10].csa.sum ;
  assign \csa0.clk  = clk;
  assign \csa0.rst  = rst;
  assign \csa0.y  = \$genblock$spm.v:14$1[1].csa.sum ;
  assign p = \csa0.sum ;
  assign pp = { \tcmp.s , \$genblock$spm.v:14$30[30].csa.sum , \$genblock$spm.v:14$29[29].csa.sum , \$genblock$spm.v:14$28[28].csa.sum , \$genblock$spm.v:14$27[27].csa.sum , \$genblock$spm.v:14$26[26].csa.sum , \$genblock$spm.v:14$25[25].csa.sum , \$genblock$spm.v:14$24[24].csa.sum , \$genblock$spm.v:14$23[23].csa.sum , \$genblock$spm.v:14$22[22].csa.sum , \$genblock$spm.v:14$21[21].csa.sum , \$genblock$spm.v:14$20[20].csa.sum , \$genblock$spm.v:14$19[19].csa.sum , \$genblock$spm.v:14$18[18].csa.sum , \$genblock$spm.v:14$17[17].csa.sum , \$genblock$spm.v:14$16[16].csa.sum , \$genblock$spm.v:14$15[15].csa.sum , \$genblock$spm.v:14$14[14].csa.sum , \$genblock$spm.v:14$13[13].csa.sum , \$genblock$spm.v:14$12[12].csa.sum , \$genblock$spm.v:14$11[11].csa.sum , \$genblock$spm.v:14$10[10].csa.sum , \$genblock$spm.v:14$9[9].csa.sum , \$genblock$spm.v:14$8[8].csa.sum , \$genblock$spm.v:14$7[7].csa.sum , \$genblock$spm.v:14$6[6].csa.sum , \$genblock$spm.v:14$5[5].csa.sum , \$genblock$spm.v:14$4[4].csa.sum , \$genblock$spm.v:14$3[3].csa.sum , \$genblock$spm.v:14$2[2].csa.sum , \$genblock$spm.v:14$1[1].csa.sum  };
  assign \tcmp.clk  = clk;
  assign \tcmp.rst  = rst;

  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


  sky130_fd_sc_hd__dlclkp
  __clk_gate_cell__
  (
    .GCLK(__clk_gate_output_GCLK_),
    .GATE(__clk_gate_input_GATE_),
    .CLK(__clk_gate_input_CLK_)
  );


endmodule

